module top() 


endmodule
